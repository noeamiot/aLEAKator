module top(input a, input b, input c, input d, output s);
    assign s = a ^ b ^ c ^ d;
endmodule
